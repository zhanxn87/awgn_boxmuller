module bm_cg_rom (clock, addr, rdata);

input              clock    ;
input  [6:0]       addr     ;
output [30:0]      rdata    ;

reg    [30:0]      rdata    ;

always @(posedge clock)
  case(addr)
    7'd0: rdata <= #1 {19'd262146, 12'd20};
    7'd1: rdata <= #1 {19'd262127, 12'd59};
    7'd2: rdata <= #1 {19'd262068, 12'd99};
    7'd3: rdata <= #1 {19'd261969, 12'd138};
    7'd4: rdata <= #1 {19'd261831, 12'd178};
    7'd5: rdata <= #1 {19'd261653, 12'd217};
    7'd6: rdata <= #1 {19'd261436, 12'd256};
    7'd7: rdata <= #1 {19'd261180, 12'd296};
    7'd8: rdata <= #1 {19'd260884, 12'd335};
    7'd9: rdata <= #1 {19'd260549, 12'd374};
    7'd10: rdata <= #1 {19'd260175, 12'd413};
    7'd11: rdata <= #1 {19'd259762, 12'd452};
    7'd12: rdata <= #1 {19'd259309, 12'd492};
    7'd13: rdata <= #1 {19'd258818, 12'd531};
    7'd14: rdata <= #1 {19'd258287, 12'd569};
    7'd15: rdata <= #1 {19'd257718, 12'd608};
    7'd16: rdata <= #1 {19'd257109, 12'd647};
    7'd17: rdata <= #1 {19'd256462, 12'd686};
    7'd18: rdata <= #1 {19'd255777, 12'd724};
    7'd19: rdata <= #1 {19'd255053, 12'd763};
    7'd20: rdata <= #1 {19'd254290, 12'd801};
    7'd21: rdata <= #1 {19'd253489, 12'd839};
    7'd22: rdata <= #1 {19'd252650, 12'd877};
    7'd23: rdata <= #1 {19'd251773, 12'd915};
    7'd24: rdata <= #1 {19'd250859, 12'd953};
    7'd25: rdata <= #1 {19'd249906, 12'd990};
    7'd26: rdata <= #1 {19'd248915, 12'd1028};
    7'd27: rdata <= #1 {19'd247888, 12'd1065};
    7'd28: rdata <= #1 {19'd246822, 12'd1102};
    7'd29: rdata <= #1 {19'd245720, 12'd1139};
    7'd30: rdata <= #1 {19'd244581, 12'd1176};
    7'd31: rdata <= #1 {19'd243405, 12'd1213};
    7'd32: rdata <= #1 {19'd242192, 12'd1249};
    7'd33: rdata <= #1 {19'd240942, 12'd1286};
    7'd34: rdata <= #1 {19'd239657, 12'd1322};
    7'd35: rdata <= #1 {19'd238335, 12'd1358};
    7'd36: rdata <= #1 {19'd236978, 12'd1393};
    7'd37: rdata <= #1 {19'd235584, 12'd1429};
    7'd38: rdata <= #1 {19'd234156, 12'd1464};
    7'd39: rdata <= #1 {19'd232692, 12'd1499};
    7'd40: rdata <= #1 {19'd231193, 12'd1534};
    7'd41: rdata <= #1 {19'd229659, 12'd1568};
    7'd42: rdata <= #1 {19'd228090, 12'd1603};
    7'd43: rdata <= #1 {19'd226487, 12'd1637};
    7'd44: rdata <= #1 {19'd224851, 12'd1671};
    7'd45: rdata <= #1 {19'd223180, 12'd1704};
    7'd46: rdata <= #1 {19'd221475, 12'd1738};
    7'd47: rdata <= #1 {19'd219738, 12'd1771};
    7'd48: rdata <= #1 {19'd217967, 12'd1804};
    7'd49: rdata <= #1 {19'd216163, 12'd1836};
    7'd50: rdata <= #1 {19'd214327, 12'd1868};
    7'd51: rdata <= #1 {19'd212458, 12'd1900};
    7'd52: rdata <= #1 {19'd210558, 12'd1932};
    7'd53: rdata <= #1 {19'd208626, 12'd1964};
    7'd54: rdata <= #1 {19'd206662, 12'd1995};
    7'd55: rdata <= #1 {19'd204668, 12'd2026};
    7'd56: rdata <= #1 {19'd202642, 12'd2056};
    7'd57: rdata <= #1 {19'd200586, 12'd2086};
    7'd58: rdata <= #1 {19'd198500, 12'd2116};
    7'd59: rdata <= #1 {19'd196383, 12'd2146};
    7'd60: rdata <= #1 {19'd194238, 12'd2175};
    7'd61: rdata <= #1 {19'd192063, 12'd2204};
    7'd62: rdata <= #1 {19'd189859, 12'd2232};
    7'd63: rdata <= #1 {19'd187626, 12'd2261};
    7'd64: rdata <= #1 {19'd185366, 12'd2289};
    7'd65: rdata <= #1 {19'd183077, 12'd2316};
    7'd66: rdata <= #1 {19'd180761, 12'd2343};
    7'd67: rdata <= #1 {19'd178417, 12'd2370};
    7'd68: rdata <= #1 {19'd176047, 12'd2397};
    7'd69: rdata <= #1 {19'd173650, 12'd2423};
    7'd70: rdata <= #1 {19'd171227, 12'd2449};
    7'd71: rdata <= #1 {19'd168778, 12'd2474};
    7'd72: rdata <= #1 {19'd166304, 12'd2499};
    7'd73: rdata <= #1 {19'd163805, 12'd2524};
    7'd74: rdata <= #1 {19'd161281, 12'd2548};
    7'd75: rdata <= #1 {19'd158733, 12'd2572};
    7'd76: rdata <= #1 {19'd156160, 12'd2596};
    7'd77: rdata <= #1 {19'd153565, 12'd2619};
    7'd78: rdata <= #1 {19'd150946, 12'd2641};
    7'd79: rdata <= #1 {19'd148305, 12'd2664};
    7'd80: rdata <= #1 {19'd145641, 12'd2686};
    7'd81: rdata <= #1 {19'd142955, 12'd2707};
    7'd82: rdata <= #1 {19'd140248, 12'd2728};
    7'd83: rdata <= #1 {19'd137519, 12'd2749};
    7'd84: rdata <= #1 {19'd134770, 12'd2769};
    7'd85: rdata <= #1 {19'd132001, 12'd2789};
    7'd86: rdata <= #1 {19'd129212, 12'd2809};
    7'd87: rdata <= #1 {19'd126403, 12'd2828};
    7'd88: rdata <= #1 {19'd123575, 12'd2846};
    7'd89: rdata <= #1 {19'd120729, 12'd2865};
    7'd90: rdata <= #1 {19'd117864, 12'd2882};
    7'd91: rdata <= #1 {19'd114982, 12'd2900};
    7'd92: rdata <= #1 {19'd112082, 12'd2917};
    7'd93: rdata <= #1 {19'd109166, 12'd2933};
    7'd94: rdata <= #1 {19'd106233, 12'd2949};
    7'd95: rdata <= #1 {19'd103284, 12'd2964};
    7'd96: rdata <= #1 {19'd100319, 12'd2980};
    7'd97: rdata <= #1 {19'd97339, 12'd2994};
    7'd98: rdata <= #1 {19'd94345, 12'd3008};
    7'd99: rdata <= #1 {19'd91337, 12'd3022};
    7'd100: rdata <= #1 {19'd88314, 12'd3036};
    7'd101: rdata <= #1 {19'd85279, 12'd3048};
    7'd102: rdata <= #1 {19'd82231, 12'd3061};
    7'd103: rdata <= #1 {19'd79170, 12'd3073};
    7'd104: rdata <= #1 {19'd76097, 12'd3084};
    7'd105: rdata <= #1 {19'd73013, 12'd3095};
    7'd106: rdata <= #1 {19'd69918, 12'd3106};
    7'd107: rdata <= #1 {19'd66812, 12'd3116};
    7'd108: rdata <= #1 {19'd63696, 12'd3125};
    7'd109: rdata <= #1 {19'd60571, 12'd3134};
    7'd110: rdata <= #1 {19'd57437, 12'd3143};
    7'd111: rdata <= #1 {19'd54294, 12'd3151};
    7'd112: rdata <= #1 {19'd51142, 12'd3159};
    7'd113: rdata <= #1 {19'd47983, 12'd3166};
    7'd114: rdata <= #1 {19'd44817, 12'd3173};
    7'd115: rdata <= #1 {19'd41644, 12'd3179};
    7'd116: rdata <= #1 {19'd38465, 12'd3185};
    7'd117: rdata <= #1 {19'd35280, 12'd3190};
    7'd118: rdata <= #1 {19'd32090, 12'd3195};
    7'd119: rdata <= #1 {19'd28894, 12'd3199};
    7'd120: rdata <= #1 {19'd25695, 12'd3203};
    7'd121: rdata <= #1 {19'd22491, 12'd3207};
    7'd122: rdata <= #1 {19'd19285, 12'd3210};
    7'd123: rdata <= #1 {19'd16075, 12'd3212};
    7'd124: rdata <= #1 {19'd12863, 12'd3214};
    7'd125: rdata <= #1 {19'd9649, 12'd3215};
    7'd126: rdata <= #1 {19'd6433, 12'd3216};
    7'd127: rdata <= #1 {19'd3217, 12'd3217};
    default: rdata <= #1 31'd0;
  endcase

endmodule

