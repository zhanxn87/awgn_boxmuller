module tb();

endmodule
