module bm_cf_rom (clock, addr, rdata);

input              clock    ;
input  [6:0]       addr     ;
output [32:0]      rdata    ;

reg    [32:0]      rdata    ;

always @(posedge clock)
  case(addr)
    7'd0: rdata <= #1 {20'd524290, 13'd4080};
    7'd1: rdata <= #1 {20'd528370, 13'd4049};
    7'd2: rdata <= #1 {20'd532419, 13'd4018};
    7'd3: rdata <= #1 {20'd536437, 13'd3988};
    7'd4: rdata <= #1 {20'd540426, 13'd3959};
    7'd5: rdata <= #1 {20'd544385, 13'd3931};
    7'd6: rdata <= #1 {20'd548315, 13'd3903};
    7'd7: rdata <= #1 {20'd552218, 13'd3875};
    7'd8: rdata <= #1 {20'd556093, 13'd3848};
    7'd9: rdata <= #1 {20'd559941, 13'd3822};
    7'd10: rdata <= #1 {20'd563764, 13'd3796};
    7'd11: rdata <= #1 {20'd567560, 13'd3771};
    7'd12: rdata <= #1 {20'd571331, 13'd3746};
    7'd13: rdata <= #1 {20'd575078, 13'd3722};
    7'd14: rdata <= #1 {20'd578800, 13'd3698};
    7'd15: rdata <= #1 {20'd582498, 13'd3675};
    7'd16: rdata <= #1 {20'd586173, 13'd3652};
    7'd17: rdata <= #1 {20'd589825, 13'd3630};
    7'd18: rdata <= #1 {20'd593455, 13'd3608};
    7'd19: rdata <= #1 {20'd597063, 13'd3586};
    7'd20: rdata <= #1 {20'd600649, 13'd3565};
    7'd21: rdata <= #1 {20'd604213, 13'd3544};
    7'd22: rdata <= #1 {20'd607757, 13'd3523};
    7'd23: rdata <= #1 {20'd611280, 13'd3503};
    7'd24: rdata <= #1 {20'd614783, 13'd3483};
    7'd25: rdata <= #1 {20'd618267, 13'd3464};
    7'd26: rdata <= #1 {20'd621730, 13'd3445};
    7'd27: rdata <= #1 {20'd625175, 13'd3426};
    7'd28: rdata <= #1 {20'd628600, 13'd3407};
    7'd29: rdata <= #1 {20'd632007, 13'd3389};
    7'd30: rdata <= #1 {20'd635396, 13'd3371};
    7'd31: rdata <= #1 {20'd638767, 13'd3353};
    7'd32: rdata <= #1 {20'd642120, 13'd3336};
    7'd33: rdata <= #1 {20'd645456, 13'd3319};
    7'd34: rdata <= #1 {20'd648774, 13'd3302};
    7'd35: rdata <= #1 {20'd652076, 13'd3285};
    7'd36: rdata <= #1 {20'd655361, 13'd3269};
    7'd37: rdata <= #1 {20'd658630, 13'd3253};
    7'd38: rdata <= #1 {20'd661882, 13'd3237};
    7'd39: rdata <= #1 {20'd665119, 13'd3221};
    7'd40: rdata <= #1 {20'd668340, 13'd3205};
    7'd41: rdata <= #1 {20'd671545, 13'd3190};
    7'd42: rdata <= #1 {20'd674735, 13'd3175};
    7'd43: rdata <= #1 {20'd677911, 13'd3160};
    7'd44: rdata <= #1 {20'd681071, 13'd3146};
    7'd45: rdata <= #1 {20'd684217, 13'd3131};
    7'd46: rdata <= #1 {20'd687348, 13'd3117};
    7'd47: rdata <= #1 {20'd690465, 13'd3103};
    7'd48: rdata <= #1 {20'd693569, 13'd3089};
    7'd49: rdata <= #1 {20'd696658, 13'd3076};
    7'd50: rdata <= #1 {20'd699734, 13'd3062};
    7'd51: rdata <= #1 {20'd702796, 13'd3049};
    7'd52: rdata <= #1 {20'd705845, 13'd3036};
    7'd53: rdata <= #1 {20'd708881, 13'd3023};
    7'd54: rdata <= #1 {20'd711904, 13'd3010};
    7'd55: rdata <= #1 {20'd714914, 13'd2998};
    7'd56: rdata <= #1 {20'd717912, 13'd2985};
    7'd57: rdata <= #1 {20'd720897, 13'd2973};
    7'd58: rdata <= #1 {20'd723870, 13'd2961};
    7'd59: rdata <= #1 {20'd726830, 13'd2949};
    7'd60: rdata <= #1 {20'd729779, 13'd2937};
    7'd61: rdata <= #1 {20'd732715, 13'd2925};
    7'd62: rdata <= #1 {20'd735640, 13'd2913};
    7'd63: rdata <= #1 {20'd738554, 13'd2902};
    7'd64: rdata <= #1 {20'd741458, 13'd5770};
    7'd65: rdata <= #1 {20'd747228, 13'd5726};
    7'd66: rdata <= #1 {20'd752954, 13'd5683};
    7'd67: rdata <= #1 {20'd758637, 13'd5640};
    7'd68: rdata <= #1 {20'd764277, 13'd5599};
    7'd69: rdata <= #1 {20'd769876, 13'd5559};
    7'd70: rdata <= #1 {20'd775435, 13'd5519};
    7'd71: rdata <= #1 {20'd780954, 13'd5480};
    7'd72: rdata <= #1 {20'd786434, 13'd5442};
    7'd73: rdata <= #1 {20'd791877, 13'd5405};
    7'd74: rdata <= #1 {20'd797282, 13'd5369};
    7'd75: rdata <= #1 {20'd802651, 13'd5333};
    7'd76: rdata <= #1 {20'd807984, 13'd5298};
    7'd77: rdata <= #1 {20'd813283, 13'd5264};
    7'd78: rdata <= #1 {20'd818546, 13'd5230};
    7'd79: rdata <= #1 {20'd823777, 13'd5197};
    7'd80: rdata <= #1 {20'd828974, 13'd5165};
    7'd81: rdata <= #1 {20'd834139, 13'd5133};
    7'd82: rdata <= #1 {20'd839272, 13'd5102};
    7'd83: rdata <= #1 {20'd844374, 13'd5071};
    7'd84: rdata <= #1 {20'd849446, 13'd5041};
    7'd85: rdata <= #1 {20'd854487, 13'd5012};
    7'd86: rdata <= #1 {20'd859498, 13'd4983};
    7'd87: rdata <= #1 {20'd864481, 13'd4954};
    7'd88: rdata <= #1 {20'd869435, 13'd4926};
    7'd89: rdata <= #1 {20'd874361, 13'd4898};
    7'd90: rdata <= #1 {20'd879259, 13'd4871};
    7'd91: rdata <= #1 {20'd884131, 13'd4845};
    7'd92: rdata <= #1 {20'd888975, 13'd4818};
    7'd93: rdata <= #1 {20'd893793, 13'd4792};
    7'd94: rdata <= #1 {20'd898586, 13'd4767};
    7'd95: rdata <= #1 {20'd903353, 13'd4742};
    7'd96: rdata <= #1 {20'd908095, 13'd4717};
    7'd97: rdata <= #1 {20'd912812, 13'd4693};
    7'd98: rdata <= #1 {20'd917505, 13'd4669};
    7'd99: rdata <= #1 {20'd922175, 13'd4646};
    7'd100: rdata <= #1 {20'd926820, 13'd4623};
    7'd101: rdata <= #1 {20'd931443, 13'd4600};
    7'd102: rdata <= #1 {20'd936043, 13'd4577};
    7'd103: rdata <= #1 {20'd940620, 13'd4555};
    7'd104: rdata <= #1 {20'd945175, 13'd4533};
    7'd105: rdata <= #1 {20'd949708, 13'd4512};
    7'd106: rdata <= #1 {20'd954220, 13'd4490};
    7'd107: rdata <= #1 {20'd958710, 13'd4470};
    7'd108: rdata <= #1 {20'd963180, 13'd4449};
    7'd109: rdata <= #1 {20'd967629, 13'd4429};
    7'd110: rdata <= #1 {20'd972057, 13'd4408};
    7'd111: rdata <= #1 {20'd976466, 13'd4389};
    7'd112: rdata <= #1 {20'd980854, 13'd4369};
    7'd113: rdata <= #1 {20'd985223, 13'd4350};
    7'd114: rdata <= #1 {20'd989573, 13'd4331};
    7'd115: rdata <= #1 {20'd993904, 13'd4312};
    7'd116: rdata <= #1 {20'd998216, 13'd4293};
    7'd117: rdata <= #1 {20'd1002509, 13'd4275};
    7'd118: rdata <= #1 {20'd1006784, 13'd4257};
    7'd119: rdata <= #1 {20'd1011041, 13'd4239};
    7'd120: rdata <= #1 {20'd1015280, 13'd4222};
    7'd121: rdata <= #1 {20'd1019502, 13'd4204};
    7'd122: rdata <= #1 {20'd1023706, 13'd4187};
    7'd123: rdata <= #1 {20'd1027893, 13'd4170};
    7'd124: rdata <= #1 {20'd1032063, 13'd4153};
    7'd125: rdata <= #1 {20'd1036216, 13'd4137};
    7'd126: rdata <= #1 {20'd1040353, 13'd4120};
    7'd127: rdata <= #1 {20'd1044473, 13'd4104};
    default: rdata <= #1 33'd0;
  endcase

endmodule

